module top();

video_ip_sim_qsys_tb tb ();
test_program pgm ();

endmodule
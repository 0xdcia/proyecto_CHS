
module unsaved (
	clk_50_in_clk,
	clk_50_2_in_clk,
	clk_50_3_in_clk,
	reset_bridge_in_reset_n);	

	input		clk_50_in_clk;
	input		clk_50_2_in_clk;
	input		clk_50_3_in_clk;
	input		reset_bridge_in_reset_n;
endmodule

// video_ip_sim_qsys_tb.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module video_ip_sim_qsys_tb (
	);

	wire    video_ip_sim_qsys_inst_clk_bfm_clk_clk;       // video_ip_sim_qsys_inst_clk_bfm:clk -> [video_ip_sim_qsys_inst:clk_clk, video_ip_sim_qsys_inst_reset_bfm:clk]
	wire    video_ip_sim_qsys_inst_reset_bfm_reset_reset; // video_ip_sim_qsys_inst_reset_bfm:reset -> video_ip_sim_qsys_inst:reset_reset_n

	video_ip_sim_qsys video_ip_sim_qsys_inst (
		.clk_clk       (video_ip_sim_qsys_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (video_ip_sim_qsys_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) video_ip_sim_qsys_inst_clk_bfm (
		.clk (video_ip_sim_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) video_ip_sim_qsys_inst_reset_bfm (
		.reset (video_ip_sim_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (video_ip_sim_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule

// video_ip_sim_qsys.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module video_ip_sim_qsys (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         video_effects_0_avalon_streaming_source_valid;             // video_effects_0:valid_out -> st_sink_bfm_0:sink_valid
	wire  [15:0] video_effects_0_avalon_streaming_source_data;              // video_effects_0:data_out -> st_sink_bfm_0:sink_data
	wire         video_effects_0_avalon_streaming_source_ready;             // st_sink_bfm_0:sink_ready -> video_effects_0:ready_in
	wire         video_effects_0_avalon_streaming_source_startofpacket;     // video_effects_0:startofpacket_out -> st_sink_bfm_0:sink_startofpacket
	wire         video_effects_0_avalon_streaming_source_endofpacket;       // video_effects_0:endofpacket_out -> st_sink_bfm_0:sink_endofpacket
	wire   [0:0] st_source_bfm_0_src_valid;                                 // st_source_bfm_0:src_valid -> video_effects_0:valid_in
	wire  [15:0] st_source_bfm_0_src_data;                                  // st_source_bfm_0:src_data -> video_effects_0:data_in
	wire         st_source_bfm_0_src_ready;                                 // video_effects_0:ready_out -> st_source_bfm_0:src_ready
	wire   [0:0] st_source_bfm_0_src_startofpacket;                         // st_source_bfm_0:src_startofpacket -> video_effects_0:startofpacket_in
	wire   [0:0] st_source_bfm_0_src_endofpacket;                           // st_source_bfm_0:src_endofpacket -> video_effects_0:endofpacket_in
	wire  [31:0] mm_master_bfm_0_m0_readdata;                               // mm_interconnect_0:mm_master_bfm_0_m0_readdata -> mm_master_bfm_0:avm_readdata
	wire         mm_master_bfm_0_m0_waitrequest;                            // mm_interconnect_0:mm_master_bfm_0_m0_waitrequest -> mm_master_bfm_0:avm_waitrequest
	wire   [2:0] mm_master_bfm_0_m0_address;                                // mm_master_bfm_0:avm_address -> mm_interconnect_0:mm_master_bfm_0_m0_address
	wire         mm_master_bfm_0_m0_read;                                   // mm_master_bfm_0:avm_read -> mm_interconnect_0:mm_master_bfm_0_m0_read
	wire  [31:0] mm_master_bfm_0_m0_writedata;                              // mm_master_bfm_0:avm_writedata -> mm_interconnect_0:mm_master_bfm_0_m0_writedata
	wire         mm_master_bfm_0_m0_write;                                  // mm_master_bfm_0:avm_write -> mm_interconnect_0:mm_master_bfm_0_m0_write
	wire         mm_interconnect_0_video_effects_0_avalon_slave_chipselect; // mm_interconnect_0:video_effects_0_avalon_slave_chipselect -> video_effects_0:chipselect
	wire  [31:0] mm_interconnect_0_video_effects_0_avalon_slave_readdata;   // video_effects_0:readdata -> mm_interconnect_0:video_effects_0_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_video_effects_0_avalon_slave_address;    // mm_interconnect_0:video_effects_0_avalon_slave_address -> video_effects_0:address
	wire         mm_interconnect_0_video_effects_0_avalon_slave_read;       // mm_interconnect_0:video_effects_0_avalon_slave_read -> video_effects_0:read
	wire         mm_interconnect_0_video_effects_0_avalon_slave_write;      // mm_interconnect_0:video_effects_0_avalon_slave_write -> video_effects_0:write
	wire  [31:0] mm_interconnect_0_video_effects_0_avalon_slave_writedata;  // mm_interconnect_0:video_effects_0_avalon_slave_writedata -> video_effects_0:writedata
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [mm_interconnect_0:mm_master_bfm_0_clk_reset_reset_bridge_in_reset_reset, mm_master_bfm_0:reset, st_sink_bfm_0:reset, st_source_bfm_0:reset, video_effects_0:reset]

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (3),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_master_bfm_0 (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.avm_address            (mm_master_bfm_0_m0_address),     //        m0.address
		.avm_readdata           (mm_master_bfm_0_m0_readdata),    //          .readdata
		.avm_writedata          (mm_master_bfm_0_m0_writedata),   //          .writedata
		.avm_waitrequest        (mm_master_bfm_0_m0_waitrequest), //          .waitrequest
		.avm_write              (mm_master_bfm_0_m0_write),       //          .write
		.avm_read               (mm_master_bfm_0_m0_read),        //          .read
		.avm_burstcount         (),                               // (terminated)
		.avm_begintransfer      (),                               // (terminated)
		.avm_beginbursttransfer (),                               // (terminated)
		.avm_byteenable         (),                               // (terminated)
		.avm_readdatavalid      (1'b0),                           // (terminated)
		.avm_arbiterlock        (),                               // (terminated)
		.avm_lock               (),                               // (terminated)
		.avm_debugaccess        (),                               // (terminated)
		.avm_transactionid      (),                               // (terminated)
		.avm_readid             (8'b00000000),                    // (terminated)
		.avm_writeid            (8'b00000000),                    // (terminated)
		.avm_clken              (),                               // (terminated)
		.avm_response           (2'b00),                          // (terminated)
		.avm_writeresponsevalid (1'b0),                           // (terminated)
		.avm_readresponse       (8'b00000000),                    // (terminated)
		.avm_writeresponse      (8'b00000000)                     // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (16),
		.ST_NUMSYMBOLS    (1),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (1),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) st_sink_bfm_0 (
		.clk                (clk_clk),                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                        // clk_reset.reset
		.sink_data          (video_effects_0_avalon_streaming_source_data),          //      sink.data
		.sink_valid         (video_effects_0_avalon_streaming_source_valid),         //          .valid
		.sink_ready         (video_effects_0_avalon_streaming_source_ready),         //          .ready
		.sink_startofpacket (video_effects_0_avalon_streaming_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_effects_0_avalon_streaming_source_endofpacket),   //          .endofpacket
		.sink_empty         (1'b0),                                                  // (terminated)
		.sink_channel       (1'b0),                                                  // (terminated)
		.sink_error         (1'b0)                                                   // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (16),
		.ST_NUMSYMBOLS    (1),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (1),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) st_source_bfm_0 (
		.clk               (clk_clk),                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),    // clk_reset.reset
		.src_data          (st_source_bfm_0_src_data),          //       src.data
		.src_valid         (st_source_bfm_0_src_valid),         //          .valid
		.src_ready         (st_source_bfm_0_src_ready),         //          .ready
		.src_startofpacket (st_source_bfm_0_src_startofpacket), //          .startofpacket
		.src_endofpacket   (st_source_bfm_0_src_endofpacket),   //          .endofpacket
		.src_empty         (),                                  // (terminated)
		.src_channel       (),                                  // (terminated)
		.src_error         ()                                   // (terminated)
	);

	video_ip video_effects_0 (
		.startofpacket_in  (st_source_bfm_0_src_startofpacket),                         //   avalon_streaming_sink.startofpacket
		.endofpacket_in    (st_source_bfm_0_src_endofpacket),                           //                        .endofpacket
		.data_in           (st_source_bfm_0_src_data),                                  //                        .data
		.ready_out         (st_source_bfm_0_src_ready),                                 //                        .ready
		.valid_in          (st_source_bfm_0_src_valid),                                 //                        .valid
		.data_out          (video_effects_0_avalon_streaming_source_data),              // avalon_streaming_source.data
		.startofpacket_out (video_effects_0_avalon_streaming_source_startofpacket),     //                        .startofpacket
		.endofpacket_out   (video_effects_0_avalon_streaming_source_endofpacket),       //                        .endofpacket
		.ready_in          (video_effects_0_avalon_streaming_source_ready),             //                        .ready
		.valid_out         (video_effects_0_avalon_streaming_source_valid),             //                        .valid
		.clk               (clk_clk),                                                   //                   clock.clk
		.reset             (rst_controller_reset_out_reset),                            //                   reset.reset
		.address           (mm_interconnect_0_video_effects_0_avalon_slave_address),    //            avalon_slave.address
		.read              (mm_interconnect_0_video_effects_0_avalon_slave_read),       //                        .read
		.readdata          (mm_interconnect_0_video_effects_0_avalon_slave_readdata),   //                        .readdata
		.write             (mm_interconnect_0_video_effects_0_avalon_slave_write),      //                        .write
		.writedata         (mm_interconnect_0_video_effects_0_avalon_slave_writedata),  //                        .writedata
		.chipselect        (mm_interconnect_0_video_effects_0_avalon_slave_chipselect)  //                        .chipselect
	);

	video_ip_sim_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                   //                                       clk_0_clk.clk
		.mm_master_bfm_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // mm_master_bfm_0_clk_reset_reset_bridge_in_reset.reset
		.mm_master_bfm_0_m0_address                            (mm_master_bfm_0_m0_address),                                //                              mm_master_bfm_0_m0.address
		.mm_master_bfm_0_m0_waitrequest                        (mm_master_bfm_0_m0_waitrequest),                            //                                                .waitrequest
		.mm_master_bfm_0_m0_read                               (mm_master_bfm_0_m0_read),                                   //                                                .read
		.mm_master_bfm_0_m0_readdata                           (mm_master_bfm_0_m0_readdata),                               //                                                .readdata
		.mm_master_bfm_0_m0_write                              (mm_master_bfm_0_m0_write),                                  //                                                .write
		.mm_master_bfm_0_m0_writedata                          (mm_master_bfm_0_m0_writedata),                              //                                                .writedata
		.video_effects_0_avalon_slave_address                  (mm_interconnect_0_video_effects_0_avalon_slave_address),    //                    video_effects_0_avalon_slave.address
		.video_effects_0_avalon_slave_write                    (mm_interconnect_0_video_effects_0_avalon_slave_write),      //                                                .write
		.video_effects_0_avalon_slave_read                     (mm_interconnect_0_video_effects_0_avalon_slave_read),       //                                                .read
		.video_effects_0_avalon_slave_readdata                 (mm_interconnect_0_video_effects_0_avalon_slave_readdata),   //                                                .readdata
		.video_effects_0_avalon_slave_writedata                (mm_interconnect_0_video_effects_0_avalon_slave_writedata),  //                                                .writedata
		.video_effects_0_avalon_slave_chipselect               (mm_interconnect_0_video_effects_0_avalon_slave_chipselect)  //                                                .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
